//==================================================
// Filename       : encoder4x2.v
// Description    : 4-to-2 Encoder (No Priority)
// GitHub         : https://github.com/AVM-27
// Author         : Adarsh Venugopal
// Created On     : 2025-08-02
//==================================================

module encoder4x2 (
    input  [3:0] in,   // One-hot input
    output reg [1:0] out // Encoded binary output
);

    always @(*) begin
        case (in)
            4'b0001: out = 2'b00;
            4'b0010: out = 2'b01;
            4'b0100: out = 2'b10;
            4'b1000: out = 2'b11;
            default: out = 2'bxx; // Invalid if not one-hot
        endcase
    end

endmodule
